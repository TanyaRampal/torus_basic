* SPICE NETLIST
***************************************

.SUBCKT LDDP D G S B
.ENDS
***************************************
.SUBCKT LDDN D G S B
.ENDS
***************************************
.SUBCKT crtmom PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT crtmom_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT crtmom_mx PLUS1 MINUS1 PLUS2 MINUS2 BULK
.ENDS
***************************************
.SUBCKT lincap PLUS MINUS
.ENDS
***************************************
.SUBCKT lincap_25 PLUS MINUS
.ENDS
***************************************
.SUBCKT lincap_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT lincap_rf_25 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT lowcpad_d0 APAD AVSS
.ENDS
***************************************
.SUBCKT lowcpad_d15 APAD AVSS
.ENDS
***************************************
.SUBCKT lowcpad_d23 APAD AVSS
.ENDS
***************************************
.SUBCKT mimcap_sin PLUS MINUS
.ENDS
***************************************
.SUBCKT mimcap_sin_3t PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_um_sin_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_woum_sin_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf18 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf18_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf25 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf25_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf33 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf33_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf_hvt PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf_hvt_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT ndio_hia_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT nmos_rf D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_18 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_18_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_18_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_25_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25_nodnwod D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25_nodnwud D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25od D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25od33_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_25ud D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25ud18_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_33 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_33_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_33_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_hvt D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_hvt_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_hvt_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_lvt D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_lvt_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_lvt_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_mlvt D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_mlvt_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_mlvt_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_na18 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmoscap PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_18 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_25 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_33 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_lpg PLUS MINUS
.ENDS
***************************************
.SUBCKT pdio_hia_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT pmos_rf D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_18 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_18_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_18_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_18_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25_nwod D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25_nwud D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25od D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25od33_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25od33_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25ud D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25ud18_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25ud18_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_33 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_33_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_33_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_33_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_hvt D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_hvt_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_hvt_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_hvt_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_lvt D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_lvt_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_lvt_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_lvt_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_mlvt D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_mlvt_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_mlvt_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_mlvt_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmoscap_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT pmoscap_rf18 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT pmoscap_rf25 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT probe1 TOP BULK
.ENDS
***************************************
.SUBCKT probe2 TOP BULK
.ENDS
***************************************
.SUBCKT probe3 TOP BULK
.ENDS
***************************************
.SUBCKT probe4 TOP BULK
.ENDS
***************************************
.SUBCKT probe5 TOP BULK
.ENDS
***************************************
.SUBCKT probe6 TOP BULK
.ENDS
***************************************
.SUBCKT probe7 TOP BULK
.ENDS
***************************************
.SUBCKT rm1 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm10 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm2 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm3 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm4 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm5 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm6 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm7 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm8 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm9 PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodl PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnods PLUS MINUS
.ENDS
***************************************
.SUBCKT rnods_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnodwo PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodwo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolyl PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolyl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolys PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolys_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolywo PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolywo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnwod PLUS MINUS
.ENDS
***************************************
.SUBCKT rnwod_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnwsti PLUS MINUS
.ENDS
***************************************
.SUBCKT rnwsti_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpodl PLUS MINUS
.ENDS
***************************************
.SUBCKT rpodl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpods PLUS MINUS
.ENDS
***************************************
.SUBCKT rpods_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpodwo PLUS MINUS
.ENDS
***************************************
.SUBCKT rpodwo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyl PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolyl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyl_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolys PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolys_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolys_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolywo PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolywo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolywo_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_rf_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_std_mu_z PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_sym_ct_mu_z PLUS MINUS BULK CTAP
.ENDS
***************************************
.SUBCKT spiral_sym_mu_z PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT xjvar PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT xjvar_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT low_swing_rx vss vdd o i
** N=5 EP=4 IP=0 FDC=4
M0 o 3 vss vss nch L=6e-08 W=3.6e-07 $X=2800 $Y=1700 $D=6
M1 vss i 3 vss nch_hvt L=6e-08 W=3.6e-07 $X=2370 $Y=1700 $D=36
M2 o 3 vdd vdd pch L=6e-08 W=7.2e-07 $X=2800 $Y=3600 $D=101
M3 vdd i 3 vdd pch_hvt L=6e-08 W=7.2e-07 $X=2370 $Y=3600 $D=113
.ENDS
***************************************
