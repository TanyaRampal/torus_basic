** Generated for: hspiceD
** Generated on: Oct 20 16:13:21 2024
** Design library name: ece720t7
** Design cell name: low_swing_tx
** Design view name: schematic
helo


.TEMP 25
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2
.LIB "/CMC/tsmc_65nm/CRN65GP/TN65CMSP018K3_V1.0C/models/hspice/crn65gplus_2d5_lk_v1d0.l" tt

** Library name: ece720t7
** Cell name: low_swing_tx
** View name: schematic
.subckt low_swing_tx c i vdd vss
m8 c net19 vss vss nch l=l4 w='w4*1' m=1 nf=1 sd=200e-9 ad='((1-int(500e-3)*2)*175e-9+(2-int(1.0)*2)*100e-9)*w4' as='((1-int(500e-3)*2)*175e-9+(2-int(1.0)*2)*250e-9)*w4' pd='(1-int(500e-3)*2)*(350e-9+2*w4)+(2-int(1.0)*2)*(200e-9+1*w4)' ps='(1-int(500e-3)*2)*(350e-9+2*w4)+(2-int(1.0)*2)*(500e-9+3*w4)' nrd='(1-int(500e-3)*2)*(100e-9/w4)+(2-int(1.0)*2)*(100e-9/w4)' nrs='(1-int(500e-3)*2)*(100e-9/w4)+(2-int(1.0)*2)*(100e-9/w4)' sa=175e-9 sb=175e-9 sca=0 scb=0 scc=0
m3 net17 net16 vss vss nch l=l1 w='w1*1' m=1 nf=1 sd=200e-9 ad='((1-int(500e-3)*2)*175e-9+(2-int(1.0)*2)*100e-9)*w1' as='((1-int(500e-3)*2)*175e-9+(2-int(1.0)*2)*250e-9)*w1' pd='(1-int(500e-3)*2)*(350e-9+2*w1)+(2-int(1.0)*2)*(200e-9+1*w1)' ps='(1-int(500e-3)*2)*(350e-9+2*w1)+(2-int(1.0)*2)*(500e-9+3*w1)' nrd='(1-int(500e-3)*2)*(100e-9/w1)+(2-int(1.0)*2)*(100e-9/w1)' nrs='(1-int(500e-3)*2)*(100e-9/w1)+(2-int(1.0)*2)*(100e-9/w1)' sa=175e-9 sb=175e-9 sca=0 scb=0 scc=0
m2 net16 net14 vss vss nch l=l2 w='w2*1' m=1 nf=1 sd=200e-9 ad='((1-int(500e-3)*2)*175e-9+(2-int(1.0)*2)*100e-9)*w2' as='((1-int(500e-3)*2)*175e-9+(2-int(1.0)*2)*250e-9)*w2' pd='(1-int(500e-3)*2)*(350e-9+2*w2)+(2-int(1.0)*2)*(200e-9+1*w2)' ps='(1-int(500e-3)*2)*(350e-9+2*w2)+(2-int(1.0)*2)*(500e-9+3*w2)' nrd='(1-int(500e-3)*2)*(100e-9/w2)+(2-int(1.0)*2)*(100e-9/w2)' nrs='(1-int(500e-3)*2)*(100e-9/w2)+(2-int(1.0)*2)*(100e-9/w2)' sa=175e-9 sb=175e-9 sca=0 scb=0 scc=0
m1 net14 net19 vss vss nch l=l2 w='w2*1' m=1 nf=1 sd=200e-9 ad='((1-int(500e-3)*2)*175e-9+(2-int(1.0)*2)*100e-9)*w2' as='((1-int(500e-3)*2)*175e-9+(2-int(1.0)*2)*250e-9)*w2' pd='(1-int(500e-3)*2)*(350e-9+2*w2)+(2-int(1.0)*2)*(200e-9+1*w2)' ps='(1-int(500e-3)*2)*(350e-9+2*w2)+(2-int(1.0)*2)*(500e-9+3*w2)' nrd='(1-int(500e-3)*2)*(100e-9/w2)+(2-int(1.0)*2)*(100e-9/w2)' nrs='(1-int(500e-3)*2)*(100e-9/w2)+(2-int(1.0)*2)*(100e-9/w2)' sa=175e-9 sb=175e-9 sca=0 scb=0 scc=0
m0 net19 i vss vss nch l=l1 w='w1*1' m=1 nf=1 sd=200e-9 ad='((1-int(500e-3)*2)*175e-9+(2-int(1.0)*2)*100e-9)*w1' as='((1-int(500e-3)*2)*175e-9+(2-int(1.0)*2)*250e-9)*w1' pd='(1-int(500e-3)*2)*(350e-9+2*w1)+(2-int(1.0)*2)*(200e-9+1*w1)' ps='(1-int(500e-3)*2)*(350e-9+2*w1)+(2-int(1.0)*2)*(500e-9+3*w1)' nrd='(1-int(500e-3)*2)*(100e-9/w1)+(2-int(1.0)*2)*(100e-9/w1)' nrs='(1-int(500e-3)*2)*(100e-9/w1)+(2-int(1.0)*2)*(100e-9/w1)' sa=175e-9 sb=175e-9 sca=0 scb=0 scc=0
m10 net33 net19 vdd vdd pch l=l3 w='w3*f' m=1 nf=f sd=200e-9 ad='((f-int(f/2)*2)*((175e-9+((f-1)*200e-9)/2)+0)+((f+1)-int((f+1)/2)*2)*((f/2)*200e-9))*w3' as='((f-int(f/2)*2)*((175e-9+((f-1)*200e-9)/2)+0)+((f+1)-int((f+1)/2)*2)*(((350e-9+(f/2-1)*200e-9)+0)+0))*w3' pd='(f-int(f/2)*2)*(((175e-9+((f-1)*200e-9)/2)+0)*2+(f+1)*w3)+((f+1)-int((f+1)/2)*2)*(((f/2)*200e-9)*2+f*w3)' ps='(f-int(f/2)*2)*(((175e-9+((f-1)*200e-9)/2)+0)*2+(f+1)*w3)+((f+1)-int((f+1)/2)*2)*((((350e-9+(f/2-1)*200e-9)+0)+0)*2+(f+2)*w3)' nrd='(f-int(f/2)*2)*((10e-15/(100e-9+100e-9*(f-1)))/w3)+((f+1)-int((f+1)/2)*2)*((100e-9/f)/w3)' nrs='(f-int(f/2)*2)*((10e-15/(100e-9+100e-9*(f-1)))/w3)+((f+1)-int((f+1)/2)*2)*((1e-21/(10e-15*(f-2)+20e-15))/w3)' sa=175e-9 sb=175e-9 sca=0 scb=0 scc=0
m9 c net17 net33 vdd pch l=l3 w='w3*f' m=1 nf=f sd=200e-9 ad='((f-int(f/2)*2)*((175e-9+((f-1)*200e-9)/2)+0)+((f+1)-int((f+1)/2)*2)*((f/2)*200e-9))*w3' as='((f-int(f/2)*2)*((175e-9+((f-1)*200e-9)/2)+0)+((f+1)-int((f+1)/2)*2)*(((350e-9+(f/2-1)*200e-9)+0)+0))*w3' pd='(f-int(f/2)*2)*(((175e-9+((f-1)*200e-9)/2)+0)*2+(f+1)*w3)+((f+1)-int((f+1)/2)*2)*(((f/2)*200e-9)*2+f*w3)' ps='(f-int(f/2)*2)*(((175e-9+((f-1)*200e-9)/2)+0)*2+(f+1)*w3)+((f+1)-int((f+1)/2)*2)*((((350e-9+(f/2-1)*200e-9)+0)+0)*2+(f+2)*w3)' nrd='(f-int(f/2)*2)*((10e-15/(100e-9+100e-9*(f-1)))/w3)+((f+1)-int((f+1)/2)*2)*((100e-9/f)/w3)' nrs='(f-int(f/2)*2)*((10e-15/(100e-9+100e-9*(f-1)))/w3)+((f+1)-int((f+1)/2)*2)*((1e-21/(10e-15*(f-2)+20e-15))/w3)' sa=175e-9 sb=175e-9 sca=0 scb=0 scc=0
m7 net17 net16 vdd vdd pch l=l1 w='(w1*2)*1' m=1 nf=1 sd=200e-9 ad='(((1-int(500e-3)*2)*175e-9+(2-int(1.0)*2)*100e-9)*w1)*2' as='(((1-int(500e-3)*2)*175e-9+(2-int(1.0)*2)*250e-9)*w1)*2' pd='(1-int(500e-3)*2)*(350e-9+(2*w1)*2)+(2-int(1.0)*2)*(200e-9+(1*w1)*2)' ps='(1-int(500e-3)*2)*(350e-9+(2*w1)*2)+(2-int(1.0)*2)*(500e-9+(3*w1)*2)' nrd='(1-int(500e-3)*2)*((100e-9/w1)*2)+(2-int(1.0)*2)*((100e-9/w1)*2)' nrs='(1-int(500e-3)*2)*((100e-9/w1)*2)+(2-int(1.0)*2)*((100e-9/w1)*2)' sa=175e-9 sb=175e-9 sca=0 scb=0 scc=0
m6 net16 net14 vdd vdd pch l=l2 w='(w2*2)*1' m=1 nf=1 sd=200e-9 ad='(((1-int(500e-3)*2)*175e-9+(2-int(1.0)*2)*100e-9)*w2)*2' as='(((1-int(500e-3)*2)*175e-9+(2-int(1.0)*2)*250e-9)*w2)*2' pd='(1-int(500e-3)*2)*(350e-9+(2*w2)*2)+(2-int(1.0)*2)*(200e-9+(1*w2)*2)' ps='(1-int(500e-3)*2)*(350e-9+(2*w2)*2)+(2-int(1.0)*2)*(500e-9+(3*w2)*2)' nrd='(1-int(500e-3)*2)*((100e-9/w2)*2)+(2-int(1.0)*2)*((100e-9/w2)*2)' nrs='(1-int(500e-3)*2)*((100e-9/w2)*2)+(2-int(1.0)*2)*((100e-9/w2)*2)' sa=175e-9 sb=175e-9 sca=0 scb=0 scc=0
m5 net14 net19 vdd vdd pch l=l2 w='(w2*2)*1' m=1 nf=1 sd=200e-9 ad='(((1-int(500e-3)*2)*175e-9+(2-int(1.0)*2)*100e-9)*w2)*2' as='(((1-int(500e-3)*2)*175e-9+(2-int(1.0)*2)*250e-9)*w2)*2' pd='(1-int(500e-3)*2)*(350e-9+(2*w2)*2)+(2-int(1.0)*2)*(200e-9+(1*w2)*2)' ps='(1-int(500e-3)*2)*(350e-9+(2*w2)*2)+(2-int(1.0)*2)*(500e-9+(3*w2)*2)' nrd='(1-int(500e-3)*2)*((100e-9/w2)*2)+(2-int(1.0)*2)*((100e-9/w2)*2)' nrs='(1-int(500e-3)*2)*((100e-9/w2)*2)+(2-int(1.0)*2)*((100e-9/w2)*2)' sa=175e-9 sb=175e-9 sca=0 scb=0 scc=0
m4 net19 i vdd vdd pch l=l1 w='(w1*2)*1' m=1 nf=1 sd=200e-9 ad='(((1-int(500e-3)*2)*175e-9+(2-int(1.0)*2)*100e-9)*w1)*2' as='(((1-int(500e-3)*2)*175e-9+(2-int(1.0)*2)*250e-9)*w1)*2' pd='(1-int(500e-3)*2)*(350e-9+(2*w1)*2)+(2-int(1.0)*2)*(200e-9+(1*w1)*2)' ps='(1-int(500e-3)*2)*(350e-9+(2*w1)*2)+(2-int(1.0)*2)*(500e-9+(3*w1)*2)' nrd='(1-int(500e-3)*2)*((100e-9/w1)*2)+(2-int(1.0)*2)*((100e-9/w1)*2)' nrs='(1-int(500e-3)*2)*((100e-9/w1)*2)+(2-int(1.0)*2)*((100e-9/w1)*2)' sa=175e-9 sb=175e-9 sca=0 scb=0 scc=0
.ends low_swing_tx
** End of subcircuit definition.
.END
